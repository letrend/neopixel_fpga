
module soc_system (
	);	

endmodule
