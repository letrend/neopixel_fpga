	component soc_system is
	end component soc_system;

	u0 : component soc_system
		port map (
		);

